module Memory(input clk, input [3:0] select, input [7:0] data_in, output reg)
